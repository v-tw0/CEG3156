library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fp_adder_top is
    port(
        data_in  : in  std_logic_vector(15 downto 0); -- Single 16-bit input
        LoadA    : in  std_logic;  -- Signal to load input to A
        LoadB    : in  std_logic;  -- Signal to load input to B
        clk      : in  std_logic;  -- Clock
        reset    : in  std_logic;  -- Reset signal
        start    : in  std_logic;  -- Start signal for addition
        done     : out std_logic;  -- Done signal
        sum      : out std_logic_vector(15 downto 0) -- Sum output
    );
end fp_adder_top;

architecture behavior of fp_adder_top is
    -- Signals for storing values
    signal A_reg, B_reg : std_logic_vector(15 downto 0);
    
    -- Component Declaration for fp_adder
    component fp_adder
        port(
            A      : in  std_logic_vector(15 downto 0);
            B      : in  std_logic_vector(15 downto 0);
            clk    : in  std_logic;
            reset  : in  std_logic;
            start  : in  std_logic;
            done   : out std_logic;
            sum    : out std_logic_vector(15 downto 0)
        );
    end component;
    
begin

    -- Instantiate the fp_adder
    uut: fp_adder port map (
        A      => A_reg,
        B      => B_reg,
        clk    => clk,
        reset  => reset,
        start  => start,
        done   => done,
        sum    => sum
    );

    -- Process to load value into A_reg or B_reg
    load_process: process(clk, reset)
    begin
        if reset = '1' then
            A_reg <= (others => '0');
            B_reg <= (others => '0');
        elsif rising_edge(clk) then
            -- Load data_in into A_reg if LoadA is enabled
            if LoadA = '1' then
                A_reg <= data_in;
            end if;
            -- Load data_in into B_reg if LoadB is enabled
            if LoadB = '1' then
                B_reg <= data_in;
            end if;
        end if;
    end process;

end behavior;
